module sinusoid
  (input [0:0] clk_i
  ,input [0:0] reset_i
   // Your ports here
   );

  // Your code here
endmodule
