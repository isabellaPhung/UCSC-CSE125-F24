module adder
  #(parameter width_p = 5)
  // You must fill in the bit widths of a_i, b_i and sum_o. a_i and
  // b_i must be width_p bits.
  (input [0:0] a_i
  ,input [0:0] b_i
  ,output [0:0] sum_o);


   // Your code here
endmodule
